// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26
module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
N870,N871,N872,N873,N875,N876,N877,
N269_1,N269_2,N269_3,N269_4,N270_1,N270_2,N270_3,N270_4,N273_1,N273_2,N273_3,N276_1,N276_2,N276_3,N279_1,N279_2,N279_3,N279_4,N280_1,N280_2,N280_3,N280_4,N284_1,N284_2,N284_3,N284_4,N286_1,N286_2,N287_1,N287_2,N287_3,N290_1,N290_2,N290_3,N291_1,N291_2,N291_3,N292_1,N292_2,N292_3,N293_1,N293_2,N293_3,N294_1,N294_2,N294_3,N295_1,N295_2,N295_3,N296_1,N296_2,N296_3,N297_1,N298_1,N302_1,N304_1,N306_1,N308_1,N309_1,N316_1,N317_1,N318_1,N323_1,N325_1,N327_1,N329_1,N331_1,N332_1,N333_1,N334_1,N335_1,N336_1,N337_1,N338_1,N339_1,N340_1,N341_1,N344_1,N349_1,N350_1,N356_1,N392_1,N400_1,N406_1,N409_1,N413_1,N416_1,N417_1,N425_1,N426_1,N427_1,N427_2,N427_3,N432_1,N432_2,N432_3,N437_1,N437_2,N442_1,N442_2,N442_3,N442_4,N443_1,N443_2,N444_1,N445_1,N475_1,N476_1,N477_1,N478_1,N479_1,N480_1,N481_1,N482_1,N488_1,N489_1,N490_1,N491_1,N499_1,N501_1,N502_1,N504_1,N506_1,N508_1,N510_1,N511_1,N512_1,N513_1,N514_1,N515_1,N516_1,N517_1,N519_1,N521_1,N522_1,N523_1,N524_1,N525_1,N526_1,N552_1,N587_1,N588_1,N589_1,N593_1,N596_1,N600_1,N605_1,N609_1,N615_1,N619_1,N624_1,N628_1,N631_1,N635_1,N640_1,N644_1,N650_1,N654_1,N659_1,N665_1,N673_1,N682_1,N692_1,N700_1,N708_1,N717_1,N727_1,N733_1,N733_2,N734_1,N734_2,N734_3,N734_4,N736_1,N737_1,N739_1,N740_1,N742_1,N743_1,N745_1,N746_1,N748_1,N749_1,N751_1,N752_1,N754_1,N755_1,N758_1,N759_1,N760_1,N763_1,N763_2,N766_1,N766_2,N773_1,N773_2,N773_3,N773_4,N778_1,N778_2,N789_1,N791_1,N793_1,N794_1,N807_1,N808_1,N809_1,N810_1,N811_1,N811_2,N811_3,N811_4,N813_1,N813_2,N814_1,N814_2,N814_3,N814_4,N815_1,N815_2,N815_3,N815_4,N819_1,N819_2,N831_1,N833_1,N835_1,N836_1,N837_1,N837_2,N838_1,N838_2,N838_3,N838_4,N839_1,N839_2,N839_3,N839_4,N849_1,N851_1,N852_1,N853_1,N854_1,N854_2,N867_1,N867_2,N868_1,N868_2,N869_1,N869_2;
nand NAND2_8 (N285, N29, N68);
nand NAND2_20 (N301, N91, N96);
nand NAND2_22 (N303, N101, N106);
nand NAND2_24 (N305, N111, N116);
nand NAND2_26 (N307, N121, N126);
not NOT1_29 (N310, N268);
nand NAND2_33 (N319, N59, N156);
nor NOR2_34 (N322, N17, N42);
nand NAND2_36 (N324, N159, N165);
nand NAND2_38 (N326, N171, N177);
nand NAND2_40 (N328, N183, N189);
nand NAND2_42 (N330, N195, N201);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
not NOT1_57 (N345, N276);
not NOT1_58 (N346, N276);
not NOT1_59 (N347, N279);
nor NOR2_60 (N348, N280, N284);
not NOT1_63 (N351, N293);
not NOT1_64 (N352, N294);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
not NOT1_73 (N369, N310);
nor NOR2_74 (N375, N322, N323);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
not NOT1_84 (N393, N345);
not NOT1_85 (N399, N346);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
nand NAND2_96 (N410, N347, N352);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
nand NAND2_128 (N466, N442, N410);
nand NAND2_137 (N483, N443, N1);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
nand NAND2_146 (N500, N463, N135);
nor NOR2_149 (N503, N475, N476);
nor NOR2_151 (N505, N477, N478);
nor NOR2_153 (N507, N479, N480);
nor NOR2_155 (N509, N481, N482);
nand NAND2_164 (N518, N130, N492);
nand NAND2_166 (N520, N495, N207);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
nor NOR2_183 (N541, N512, N513);
nor NOR2_184 (N542, N514, N515);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
nand NAND2_197 (N577, N490, N542);
nand NAND2_198 (N581, N491, N543);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
nand NAND2_204 (N590, N553, N159);
nand NAND2_207 (N597, N557, N165);
nand NAND2_210 (N606, N561, N171);
nand NAND2_213 (N616, N565, N177);
nand NAND2_216 (N625, N569, N183);
nand NAND2_219 (N632, N573, N189);
nand NAND2_222 (N641, N577, N195);
nand NAND2_225 (N651, N581, N201);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
not NOT1_257 (N735, N662);
not NOT1_260 (N738, N670);
not NOT1_263 (N741, N678);
not NOT1_266 (N744, N687);
not NOT1_269 (N747, N697);
not NOT1_272 (N750, N705);
not NOT1_275 (N753, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
nand NAND2_283 (N761, N644, N722);
nand NAND2_284 (N762, N635, N713);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
nor NOR2_296 (N777, N748, N749);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700, N773);
nor NOR2_305 (N790, N708, N778);
nor NOR2_307 (N792, N717, N782);
nand NAND2_310 (N795, N628, N773);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692, N796);
nand NAND2_322 (N812, N619, N796);
nand NAND2_327 (N822, N744, N812);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
nor NOR2_333 (N830, N665, N815);
nor NOR2_335 (N832, N673, N819);
nor NOR2_337 (N834, N682, N822);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815, N593);
nor NOR2_345 (N842, N830, N831);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
buf BUFF1_353 (N850, N840);
not NOT1_358 (N855, N846);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
not NOT1_361 (N858, N849);
nor NOR2_362 (N859, N417, N851);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
not NOT1_373 (N870, N862);
not NOT1_374 (N871, N867);
not NOT1_375 (N872, N868);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);
not NOT1_NEW_3 (N269_3, N269_1);
not NOT1_NEW_4 (N269_4, N269_2);
nand NAND2_NEW_1 (N269_1, N1, N8);
nand NAND2_NEW_2 (N269_2, N13, N17);
nand NAND2_NEW_5 (N269, N269_3, N269_4);
not NOT1_NEW_8 (N270_3, N270_1);
not NOT1_NEW_9 (N270_4, N270_2);
nand NAND2_NEW_6 (N270_1, N1, N26);
nand NAND2_NEW_7 (N270_2, N13, N17);
nand NAND2_NEW_10 (N270, N270_3, N270_4);
not NOT1_NEW_12 (N273_2, N273_1);
not NOT1_NEW_14 (N273, N273_3);
nand NAND2_NEW_11 (N273_1, N29, N36);
nand NAND2_NEW_13 (N273_3, N42, N273_2);
not NOT1_NEW_16 (N276_2, N276_1);
not NOT1_NEW_18 (N276, N276_3);
nand NAND2_NEW_15 (N276_1, N1, N26);
nand NAND2_NEW_17 (N276_3, N51, N276_2);
not NOT1_NEW_21 (N279_3, N279_1);
not NOT1_NEW_22 (N279_4, N279_2);
nand NAND2_NEW_19 (N279_1, N1, N8);
nand NAND2_NEW_20 (N279_2, N51, N17);
nand NAND2_NEW_23 (N279, N279_3, N279_4);
not NOT1_NEW_26 (N280_3, N280_1);
not NOT1_NEW_27 (N280_4, N280_2);
nand NAND2_NEW_24 (N280_1, N1, N8);
nand NAND2_NEW_25 (N280_2, N13, N55);
nand NAND2_NEW_28 (N280, N280_3, N280_4);
not NOT1_NEW_31 (N284_3, N284_1);
not NOT1_NEW_32 (N284_4, N284_2);
nand NAND2_NEW_29 (N284_1, N59, N42);
nand NAND2_NEW_30 (N284_2, N68, N72);
nand NAND2_NEW_33 (N284, N284_3, N284_4);
not NOT1_NEW_35 (N286_2, N286_1);
nand NAND2_NEW_34 (N286_1, N59, N68);
nand NAND2_NEW_36 (N286, N74, N286_2);
not NOT1_NEW_38 (N287_2, N287_1);
not NOT1_NEW_40 (N287, N287_3);
nand NAND2_NEW_37 (N287_1, N29, N75);
nand NAND2_NEW_39 (N287_3, N80, N287_2);
not NOT1_NEW_42 (N290_2, N290_1);
not NOT1_NEW_44 (N290, N290_3);
nand NAND2_NEW_41 (N290_1, N29, N75);
nand NAND2_NEW_43 (N290_3, N42, N290_2);
not NOT1_NEW_46 (N291_2, N291_1);
not NOT1_NEW_48 (N291, N291_3);
nand NAND2_NEW_45 (N291_1, N29, N36);
nand NAND2_NEW_47 (N291_3, N80, N291_2);
not NOT1_NEW_50 (N292_2, N292_1);
not NOT1_NEW_52 (N292, N292_3);
nand NAND2_NEW_49 (N292_1, N29, N36);
nand NAND2_NEW_51 (N292_3, N42, N292_2);
not NOT1_NEW_54 (N293_2, N293_1);
not NOT1_NEW_56 (N293, N293_3);
nand NAND2_NEW_53 (N293_1, N59, N75);
nand NAND2_NEW_55 (N293_3, N80, N293_2);
not NOT1_NEW_58 (N294_2, N294_1);
not NOT1_NEW_60 (N294, N294_3);
nand NAND2_NEW_57 (N294_1, N59, N75);
nand NAND2_NEW_59 (N294_3, N42, N294_2);
not NOT1_NEW_62 (N295_2, N295_1);
not NOT1_NEW_64 (N295, N295_3);
nand NAND2_NEW_61 (N295_1, N59, N36);
nand NAND2_NEW_63 (N295_3, N80, N295_2);
not NOT1_NEW_66 (N296_2, N296_1);
not NOT1_NEW_68 (N296, N296_3);
nand NAND2_NEW_65 (N296_1, N59, N36);
nand NAND2_NEW_67 (N296_3, N42, N296_2);
nand NAND2_NEW_69 (N297_1, N85, N86);
not NOT1_NEW_70 (N297, N297_1);
nor NOR2_NEW_71 (N298_1, N87, N88);
not NOT1_NEW_72 (N298, N298_1);
nor NOR2_NEW_73 (N302_1, N91, N96);
not NOT1_NEW_74 (N302, N302_1);
nor NOR2_NEW_75 (N304_1, N101, N106);
not NOT1_NEW_76 (N304, N304_1);
nor NOR2_NEW_77 (N306_1, N111, N116);
not NOT1_NEW_78 (N306, N306_1);
nor NOR2_NEW_79 (N308_1, N121, N126);
not NOT1_NEW_80 (N308, N308_1);
nand NAND2_NEW_81 (N309_1, N8, N138);
not NOT1_NEW_82 (N309, N309_1);
nand NAND2_NEW_83 (N316_1, N51, N138);
not NOT1_NEW_84 (N316, N316_1);
nand NAND2_NEW_85 (N317_1, N17, N138);
not NOT1_NEW_86 (N317, N317_1);
nand NAND2_NEW_87 (N318_1, N152, N138);
not NOT1_NEW_88 (N318, N318_1);
nand NAND2_NEW_89 (N323_1, N17, N42);
not NOT1_NEW_90 (N323, N323_1);
nor NOR2_NEW_91 (N325_1, N159, N165);
not NOT1_NEW_92 (N325, N325_1);
nor NOR2_NEW_93 (N327_1, N171, N177);
not NOT1_NEW_94 (N327, N327_1);
nor NOR2_NEW_95 (N329_1, N183, N189);
not NOT1_NEW_96 (N329, N329_1);
nor NOR2_NEW_97 (N331_1, N195, N201);
not NOT1_NEW_98 (N331, N331_1);
nand NAND2_NEW_99 (N332_1, N210, N91);
not NOT1_NEW_100 (N332, N332_1);
nand NAND2_NEW_101 (N333_1, N210, N96);
not NOT1_NEW_102 (N333, N333_1);
nand NAND2_NEW_103 (N334_1, N210, N101);
not NOT1_NEW_104 (N334, N334_1);
nand NAND2_NEW_105 (N335_1, N210, N106);
not NOT1_NEW_106 (N335, N335_1);
nand NAND2_NEW_107 (N336_1, N210, N111);
not NOT1_NEW_108 (N336, N336_1);
nand NAND2_NEW_109 (N337_1, N255, N259);
not NOT1_NEW_110 (N337, N337_1);
nand NAND2_NEW_111 (N338_1, N210, N116);
not NOT1_NEW_112 (N338, N338_1);
nand NAND2_NEW_113 (N339_1, N255, N260);
not NOT1_NEW_114 (N339, N339_1);
nand NAND2_NEW_115 (N340_1, N210, N121);
not NOT1_NEW_116 (N340, N340_1);
nand NAND2_NEW_117 (N341_1, N255, N267);
not NOT1_NEW_118 (N341, N341_1);
nor NOR2_NEW_119 (N344_1, N270, N273);
not NOT1_NEW_120 (N344, N344_1);
nor NOR2_NEW_121 (N349_1, N280, N285);
not NOT1_NEW_122 (N349, N349_1);
nor NOR2_NEW_123 (N350_1, N280, N286);
not NOT1_NEW_124 (N350, N350_1);
nand NAND2_NEW_125 (N356_1, N90, N298);
not NOT1_NEW_126 (N356, N356_1);
nor NOR2_NEW_127 (N392_1, N270, N343);
not NOT1_NEW_128 (N392, N392_1);
nand NAND2_NEW_129 (N400_1, N348, N73);
not NOT1_NEW_130 (N400, N400_1);
nand NAND2_NEW_131 (N406_1, N357, N360);
not NOT1_NEW_132 (N406, N406_1);
nand NAND2_NEW_133 (N409_1, N363, N366);
not NOT1_NEW_134 (N409, N409_1);
nand NAND2_NEW_135 (N413_1, N376, N379);
not NOT1_NEW_136 (N413, N413_1);
nand NAND2_NEW_137 (N416_1, N382, N385);
not NOT1_NEW_138 (N416, N416_1);
nand NAND2_NEW_139 (N417_1, N210, N369);
not NOT1_NEW_140 (N417, N417_1);
nand NAND2_NEW_141 (N425_1, N404, N405);
not NOT1_NEW_142 (N425, N425_1);
nand NAND2_NEW_143 (N426_1, N407, N408);
not NOT1_NEW_144 (N426, N426_1);
not NOT1_NEW_146 (N427_2, N427_1);
not NOT1_NEW_148 (N427, N427_3);
nand NAND2_NEW_145 (N427_1, N319, N393);
nand NAND2_NEW_147 (N427_3, N55, N427_2);
not NOT1_NEW_150 (N432_2, N432_1);
not NOT1_NEW_152 (N432, N432_3);
nand NAND2_NEW_149 (N432_1, N393, N17);
nand NAND2_NEW_151 (N432_3, N287, N432_2);
not NOT1_NEW_154 (N437_2, N437_1);
nand NAND2_NEW_153 (N437_1, N393, N287);
nand NAND2_NEW_155 (N437, N55, N437_2);
not NOT1_NEW_158 (N442_3, N442_1);
not NOT1_NEW_159 (N442_4, N442_2);
nand NAND2_NEW_156 (N442_1, N375, N59);
nand NAND2_NEW_157 (N442_2, N156, N393);
nand NAND2_NEW_160 (N442, N442_3, N442_4);
not NOT1_NEW_162 (N443_2, N443_1);
nand NAND2_NEW_161 (N443_1, N393, N319);
nand NAND2_NEW_163 (N443, N17, N443_2);
nand NAND2_NEW_164 (N444_1, N411, N412);
not NOT1_NEW_165 (N444, N444_1);
nand NAND2_NEW_166 (N445_1, N414, N415);
not NOT1_NEW_167 (N445, N445_1);
nand NAND2_NEW_168 (N475_1, N143, N427);
not NOT1_NEW_169 (N475, N475_1);
nand NAND2_NEW_170 (N476_1, N310, N432);
not NOT1_NEW_171 (N476, N476_1);
nand NAND2_NEW_172 (N477_1, N146, N427);
not NOT1_NEW_173 (N477, N477_1);
nand NAND2_NEW_174 (N478_1, N310, N432);
not NOT1_NEW_175 (N478, N478_1);
nand NAND2_NEW_176 (N479_1, N149, N427);
not NOT1_NEW_177 (N479, N479_1);
nand NAND2_NEW_178 (N480_1, N310, N432);
not NOT1_NEW_179 (N480, N480_1);
nand NAND2_NEW_180 (N481_1, N153, N427);
not NOT1_NEW_181 (N481, N481_1);
nand NAND2_NEW_182 (N482_1, N310, N432);
not NOT1_NEW_183 (N482, N482_1);
nor NOR2_NEW_184 (N488_1, N369, N437);
not NOT1_NEW_185 (N488, N488_1);
nor NOR2_NEW_186 (N489_1, N369, N437);
not NOT1_NEW_187 (N489, N489_1);
nor NOR2_NEW_188 (N490_1, N369, N437);
not NOT1_NEW_189 (N490, N490_1);
nor NOR2_NEW_190 (N491_1, N369, N437);
not NOT1_NEW_191 (N491, N491_1);
nor NOR2_NEW_192 (N499_1, N130, N460);
not NOT1_NEW_193 (N499, N499_1);
nor NOR2_NEW_194 (N501_1, N463, N135);
not NOT1_NEW_195 (N501, N501_1);
nand NAND2_NEW_196 (N502_1, N91, N466);
not NOT1_NEW_197 (N502, N502_1);
nand NAND2_NEW_198 (N504_1, N96, N466);
not NOT1_NEW_199 (N504, N504_1);
nand NAND2_NEW_200 (N506_1, N101, N466);
not NOT1_NEW_201 (N506, N506_1);
nand NAND2_NEW_202 (N508_1, N106, N466);
not NOT1_NEW_203 (N508, N508_1);
nand NAND2_NEW_204 (N510_1, N143, N483);
not NOT1_NEW_205 (N510, N510_1);
nand NAND2_NEW_206 (N511_1, N111, N466);
not NOT1_NEW_207 (N511, N511_1);
nand NAND2_NEW_208 (N512_1, N146, N483);
not NOT1_NEW_209 (N512, N512_1);
nand NAND2_NEW_210 (N513_1, N116, N466);
not NOT1_NEW_211 (N513, N513_1);
nand NAND2_NEW_212 (N514_1, N149, N483);
not NOT1_NEW_213 (N514, N514_1);
nand NAND2_NEW_214 (N515_1, N121, N466);
not NOT1_NEW_215 (N515, N515_1);
nand NAND2_NEW_216 (N516_1, N153, N483);
not NOT1_NEW_217 (N516, N516_1);
nand NAND2_NEW_218 (N517_1, N126, N466);
not NOT1_NEW_219 (N517, N517_1);
nor NOR2_NEW_220 (N519_1, N130, N492);
not NOT1_NEW_221 (N519, N519_1);
nor NOR2_NEW_222 (N521_1, N495, N207);
not NOT1_NEW_223 (N521, N521_1);
nand NAND2_NEW_224 (N522_1, N451, N159);
not NOT1_NEW_225 (N522, N522_1);
nand NAND2_NEW_226 (N523_1, N451, N165);
not NOT1_NEW_227 (N523, N523_1);
nand NAND2_NEW_228 (N524_1, N451, N171);
not NOT1_NEW_229 (N524, N524_1);
nand NAND2_NEW_230 (N525_1, N451, N177);
not NOT1_NEW_231 (N525, N525_1);
nand NAND2_NEW_232 (N526_1, N451, N183);
not NOT1_NEW_233 (N526, N526_1);
nand NAND2_NEW_234 (N552_1, N530, N533);
not NOT1_NEW_235 (N552, N552_1);
nand NAND2_NEW_236 (N587_1, N544, N547);
not NOT1_NEW_237 (N587, N587_1);
nand NAND2_NEW_238 (N588_1, N550, N551);
not NOT1_NEW_239 (N588, N588_1);
nand NAND2_NEW_240 (N589_1, N585, N586);
not NOT1_NEW_241 (N589, N589_1);
nor NOR2_NEW_242 (N593_1, N553, N159);
not NOT1_NEW_243 (N593, N593_1);
nand NAND2_NEW_244 (N596_1, N246, N553);
not NOT1_NEW_245 (N596, N596_1);
nor NOR2_NEW_246 (N600_1, N557, N165);
not NOT1_NEW_247 (N600, N600_1);
nand NAND2_NEW_248 (N605_1, N246, N557);
not NOT1_NEW_249 (N605, N605_1);
nor NOR2_NEW_250 (N609_1, N561, N171);
not NOT1_NEW_251 (N609, N609_1);
nand NAND2_NEW_252 (N615_1, N246, N561);
not NOT1_NEW_253 (N615, N615_1);
nor NOR2_NEW_254 (N619_1, N565, N177);
not NOT1_NEW_255 (N619, N619_1);
nand NAND2_NEW_256 (N624_1, N246, N565);
not NOT1_NEW_257 (N624, N624_1);
nor NOR2_NEW_258 (N628_1, N569, N183);
not NOT1_NEW_259 (N628, N628_1);
nand NAND2_NEW_260 (N631_1, N246, N569);
not NOT1_NEW_261 (N631, N631_1);
nor NOR2_NEW_262 (N635_1, N573, N189);
not NOT1_NEW_263 (N635, N635_1);
nand NAND2_NEW_264 (N640_1, N246, N573);
not NOT1_NEW_265 (N640, N640_1);
nor NOR2_NEW_266 (N644_1, N577, N195);
not NOT1_NEW_267 (N644, N644_1);
nand NAND2_NEW_268 (N650_1, N246, N577);
not NOT1_NEW_269 (N650, N650_1);
nor NOR2_NEW_270 (N654_1, N581, N201);
not NOT1_NEW_271 (N654, N654_1);
nand NAND2_NEW_272 (N659_1, N246, N581);
not NOT1_NEW_273 (N659, N659_1);
nand NAND2_NEW_274 (N665_1, N593, N590);
not NOT1_NEW_275 (N665, N665_1);
nand NAND2_NEW_276 (N673_1, N600, N597);
not NOT1_NEW_277 (N673, N673_1);
nand NAND2_NEW_278 (N682_1, N609, N606);
not NOT1_NEW_279 (N682, N682_1);
nand NAND2_NEW_280 (N692_1, N619, N616);
not NOT1_NEW_281 (N692, N692_1);
nand NAND2_NEW_282 (N700_1, N628, N625);
not NOT1_NEW_283 (N700, N700_1);
nand NAND2_NEW_284 (N708_1, N635, N632);
not NOT1_NEW_285 (N708, N708_1);
nand NAND2_NEW_286 (N717_1, N644, N641);
not NOT1_NEW_287 (N717, N717_1);
nand NAND2_NEW_288 (N727_1, N654, N651);
not NOT1_NEW_289 (N727, N727_1);
not NOT1_NEW_291 (N733_2, N733_1);
nand NAND2_NEW_290 (N733_1, N644, N654);
nand NAND2_NEW_292 (N733, N261, N733_2);
not NOT1_NEW_295 (N734_3, N734_1);
not NOT1_NEW_296 (N734_4, N734_2);
nand NAND2_NEW_293 (N734_1, N635, N644);
nand NAND2_NEW_294 (N734_2, N654, N261);
nand NAND2_NEW_297 (N734, N734_3, N734_4);
nand NAND2_NEW_298 (N736_1, N228, N665);
not NOT1_NEW_299 (N736, N736_1);
nand NAND2_NEW_300 (N737_1, N237, N662);
not NOT1_NEW_301 (N737, N737_1);
nand NAND2_NEW_302 (N739_1, N228, N673);
not NOT1_NEW_303 (N739, N739_1);
nand NAND2_NEW_304 (N740_1, N237, N670);
not NOT1_NEW_305 (N740, N740_1);
nand NAND2_NEW_306 (N742_1, N228, N682);
not NOT1_NEW_307 (N742, N742_1);
nand NAND2_NEW_308 (N743_1, N237, N678);
not NOT1_NEW_309 (N743, N743_1);
nand NAND2_NEW_310 (N745_1, N228, N692);
not NOT1_NEW_311 (N745, N745_1);
nand NAND2_NEW_312 (N746_1, N237, N687);
not NOT1_NEW_313 (N746, N746_1);
nand NAND2_NEW_314 (N748_1, N228, N700);
not NOT1_NEW_315 (N748, N748_1);
nand NAND2_NEW_316 (N749_1, N237, N697);
not NOT1_NEW_317 (N749, N749_1);
nand NAND2_NEW_318 (N751_1, N228, N708);
not NOT1_NEW_319 (N751, N751_1);
nand NAND2_NEW_320 (N752_1, N237, N705);
not NOT1_NEW_321 (N752, N752_1);
nand NAND2_NEW_322 (N754_1, N228, N717);
not NOT1_NEW_323 (N754, N754_1);
nand NAND2_NEW_324 (N755_1, N237, N713);
not NOT1_NEW_325 (N755, N755_1);
nand NAND2_NEW_326 (N758_1, N727, N261);
not NOT1_NEW_327 (N758, N758_1);
nand NAND2_NEW_328 (N759_1, N228, N727);
not NOT1_NEW_329 (N759, N759_1);
nand NAND2_NEW_330 (N760_1, N237, N722);
not NOT1_NEW_331 (N760, N760_1);
not NOT1_NEW_333 (N763_2, N763_1);
nand NAND2_NEW_332 (N763_1, N635, N644);
nand NAND2_NEW_334 (N763, N722, N763_2);
not NOT1_NEW_336 (N766_2, N766_1);
nand NAND2_NEW_335 (N766_1, N600, N609);
nand NAND2_NEW_337 (N766, N687, N766_2);
not NOT1_NEW_340 (N773_3, N773_1);
not NOT1_NEW_341 (N773_4, N773_2);
nand NAND2_NEW_338 (N773_1, N750, N762);
nand NAND2_NEW_339 (N773_2, N763, N734);
nand NAND2_NEW_342 (N773, N773_3, N773_4);
not NOT1_NEW_344 (N778_2, N778_1);
nand NAND2_NEW_343 (N778_1, N753, N761);
nand NAND2_NEW_345 (N778, N733, N778_2);
nand NAND2_NEW_346 (N789_1, N700, N773);
not NOT1_NEW_347 (N789, N789_1);
nand NAND2_NEW_348 (N791_1, N708, N778);
not NOT1_NEW_349 (N791, N791_1);
nand NAND2_NEW_350 (N793_1, N717, N782);
not NOT1_NEW_351 (N793, N793_1);
nand NAND2_NEW_352 (N794_1, N219, N786);
not NOT1_NEW_353 (N794, N794_1);
nand NAND2_NEW_354 (N807_1, N692, N796);
not NOT1_NEW_355 (N807, N807_1);
nand NAND2_NEW_356 (N808_1, N219, N802);
not NOT1_NEW_357 (N808, N808_1);
nand NAND2_NEW_358 (N809_1, N219, N803);
not NOT1_NEW_359 (N809, N809_1);
nand NAND2_NEW_360 (N810_1, N219, N804);
not NOT1_NEW_361 (N810, N810_1);
not NOT1_NEW_364 (N811_3, N811_1);
not NOT1_NEW_365 (N811_4, N811_2);
nand NAND2_NEW_362 (N811_1, N805, N787);
nand NAND2_NEW_363 (N811_2, N731, N529);
nand NAND2_NEW_366 (N811, N811_3, N811_4);
not NOT1_NEW_368 (N813_2, N813_1);
nand NAND2_NEW_367 (N813_1, N609, N619);
nand NAND2_NEW_369 (N813, N796, N813_2);
not NOT1_NEW_372 (N814_3, N814_1);
not NOT1_NEW_373 (N814_4, N814_2);
nand NAND2_NEW_370 (N814_1, N600, N609);
nand NAND2_NEW_371 (N814_2, N619, N796);
nand NAND2_NEW_374 (N814, N814_3, N814_4);
not NOT1_NEW_377 (N815_3, N815_1);
not NOT1_NEW_378 (N815_4, N815_2);
nand NAND2_NEW_375 (N815_1, N738, N765);
nand NAND2_NEW_376 (N815_2, N766, N814);
nand NAND2_NEW_379 (N815, N815_3, N815_4);
not NOT1_NEW_381 (N819_2, N819_1);
nand NAND2_NEW_380 (N819_1, N741, N764);
nand NAND2_NEW_382 (N819, N813, N819_2);
nand NAND2_NEW_383 (N831_1, N665, N815);
not NOT1_NEW_384 (N831, N831_1);
nand NAND2_NEW_385 (N833_1, N673, N819);
not NOT1_NEW_386 (N833, N833_1);
nand NAND2_NEW_387 (N835_1, N682, N822);
not NOT1_NEW_388 (N835, N835_1);
nand NAND2_NEW_389 (N836_1, N219, N825);
not NOT1_NEW_390 (N836, N836_1);
not NOT1_NEW_392 (N837_2, N837_1);
nand NAND2_NEW_391 (N837_1, N826, N777);
nand NAND2_NEW_393 (N837, N704, N837_2);
not NOT1_NEW_396 (N838_3, N838_1);
not NOT1_NEW_397 (N838_4, N838_2);
nand NAND2_NEW_394 (N838_1, N827, N781);
nand NAND2_NEW_395 (N838_2, N712, N527);
nand NAND2_NEW_398 (N838, N838_3, N838_4);
not NOT1_NEW_401 (N839_3, N839_1);
not NOT1_NEW_402 (N839_4, N839_2);
nand NAND2_NEW_399 (N839_1, N828, N785);
nand NAND2_NEW_400 (N839_2, N721, N528);
nand NAND2_NEW_403 (N839, N839_3, N839_4);
nand NAND2_NEW_404 (N849_1, N735, N841);
not NOT1_NEW_405 (N849, N849_1);
nand NAND2_NEW_406 (N851_1, N219, N842);
not NOT1_NEW_407 (N851, N851_1);
nand NAND2_NEW_408 (N852_1, N219, N843);
not NOT1_NEW_409 (N852, N852_1);
nand NAND2_NEW_410 (N853_1, N219, N844);
not NOT1_NEW_411 (N853, N853_1);
not NOT1_NEW_413 (N854_2, N854_1);
nand NAND2_NEW_412 (N854_1, N845, N772);
nand NAND2_NEW_414 (N854, N696, N854_2);
not NOT1_NEW_416 (N867_2, N867_1);
nand NAND2_NEW_415 (N867_1, N859, N769);
nand NAND2_NEW_417 (N867, N669, N867_2);
not NOT1_NEW_419 (N868_2, N868_1);
nand NAND2_NEW_418 (N868_1, N860, N770);
nand NAND2_NEW_420 (N868, N677, N868_2);
not NOT1_NEW_422 (N869_2, N869_1);
nand NAND2_NEW_421 (N869_1, N861, N771);
nand NAND2_NEW_423 (N869, N686, N869_2);
endmodule
