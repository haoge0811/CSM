// Verilog
// inv
// Ninputs 1
// Noutputs 1
// NtotalGates 1
// NOT 1

module inv (N1,N2);

input N1;

output N2;

not NOT1_1 (N2, N1);

endmodule